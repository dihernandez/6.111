`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// camera module
//////////////////////////////////////////////////////////////////////////////////

module camera (
        input clk,
        input data_in,
        output logic [7:0] data_out
    );

    assign data_out = 8'b0;

endmodule
